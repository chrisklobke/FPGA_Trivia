-- finalproject_trivia.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity finalproject_trivia is
	port (
		clk_clk                                      : in    std_logic                     := '0';             --                                   clk.clk
		clk_sdram_clk                                : out   std_logic;                                        --                             clk_sdram.clk
		pio_input_key_external_connection_export     : in    std_logic_vector(3 downto 0)  := (others => '0'); --     pio_input_key_external_connection.export
		pio_input_level_external_connection_export   : in    std_logic_vector(3 downto 0)  := (others => '0'); --   pio_input_level_external_connection.export
		pio_output_answer_external_connection_export : out   std_logic_vector(1 downto 0);                     -- pio_output_answer_external_connection.export
		pio_sseg_external_connection_export          : out   std_logic_vector(15 downto 0);                    --          pio_sseg_external_connection.export
		reset_reset_n                                : in    std_logic                     := '0';             --                                 reset.reset_n
		sdram_wire_addr                              : out   std_logic_vector(12 downto 0);                    --                            sdram_wire.addr
		sdram_wire_ba                                : out   std_logic_vector(1 downto 0);                     --                                      .ba
		sdram_wire_cas_n                             : out   std_logic;                                        --                                      .cas_n
		sdram_wire_cke                               : out   std_logic;                                        --                                      .cke
		sdram_wire_cs_n                              : out   std_logic;                                        --                                      .cs_n
		sdram_wire_dq                                : inout std_logic_vector(15 downto 0) := (others => '0'); --                                      .dq
		sdram_wire_dqm                               : out   std_logic_vector(1 downto 0);                     --                                      .dqm
		sdram_wire_ras_n                             : out   std_logic;                                        --                                      .ras_n
		sdram_wire_we_n                              : out   std_logic;                                        --                                      .we_n
		vga_out_CLK                                  : out   std_logic;                                        --                               vga_out.CLK
		vga_out_HS                                   : out   std_logic;                                        --                                      .HS
		vga_out_VS                                   : out   std_logic;                                        --                                      .VS
		vga_out_BLANK                                : out   std_logic;                                        --                                      .BLANK
		vga_out_SYNC                                 : out   std_logic;                                        --                                      .SYNC
		vga_out_R                                    : out   std_logic_vector(3 downto 0);                     --                                      .R
		vga_out_G                                    : out   std_logic_vector(3 downto 0);                     --                                      .G
		vga_out_B                                    : out   std_logic_vector(3 downto 0)                      --                                      .B
	);
end entity finalproject_trivia;

architecture rtl of finalproject_trivia is
	component finalproject_trivia_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component finalproject_trivia_altpll_0;

	component finalproject_trivia_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component finalproject_trivia_jtag_uart_0;

	component finalproject_trivia_new_sdram_controller_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component finalproject_trivia_new_sdram_controller_0;

	component finalproject_trivia_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(26 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component finalproject_trivia_nios2_gen2_0;

	component finalproject_trivia_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component finalproject_trivia_onchip_memory2_0;

	component finalproject_trivia_pio_input_key is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component finalproject_trivia_pio_input_key;

	component finalproject_trivia_pio_output_answer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component finalproject_trivia_pio_output_answer;

	component finalproject_trivia_pio_sseg is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component finalproject_trivia_pio_sseg;

	component finalproject_trivia_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component finalproject_trivia_sysid_qsys_0;

	component finalproject_trivia_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component finalproject_trivia_timer_0;

	component finalproject_trivia_video_character_buffer_with_dma_0 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			ctrl_address         : in  std_logic                     := 'X';             -- address
			ctrl_byteenable      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ctrl_chipselect      : in  std_logic                     := 'X';             -- chipselect
			ctrl_read            : in  std_logic                     := 'X';             -- read
			ctrl_write           : in  std_logic                     := 'X';             -- write
			ctrl_writedata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ctrl_readdata        : out std_logic_vector(31 downto 0);                    -- readdata
			buf_byteenable       : in  std_logic                     := 'X';             -- byteenable
			buf_chipselect       : in  std_logic                     := 'X';             -- chipselect
			buf_read             : in  std_logic                     := 'X';             -- read
			buf_write            : in  std_logic                     := 'X';             -- write
			buf_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			buf_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			buf_waitrequest      : out std_logic;                                        -- waitrequest
			buf_address          : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component finalproject_trivia_video_character_buffer_with_dma_0;

	component finalproject_trivia_video_dual_clock_buffer_0 is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component finalproject_trivia_video_dual_clock_buffer_0;

	component finalproject_trivia_video_vga_controller_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(3 downto 0);                     -- export
			VGA_G         : out std_logic_vector(3 downto 0);                     -- export
			VGA_B         : out std_logic_vector(3 downto 0)                      -- export
		);
	end component finalproject_trivia_video_vga_controller_0;

	component finalproject_trivia_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                                        : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                                          : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset             : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                         : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                                       : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                                   : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                                    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                                          : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                                      : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                                         : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                                   : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address                                : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest                            : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                                   : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata                               : out std_logic_vector(31 downto 0);                    -- readdata
			altpll_0_pll_slave_address                                             : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                               : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                                : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_address                                  : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                                    : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                                     : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                              : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                               : out std_logic;                                        -- chipselect
			new_sdram_controller_0_s1_address                                      : out std_logic_vector(24 downto 0);                    -- address
			new_sdram_controller_0_s1_write                                        : out std_logic;                                        -- write
			new_sdram_controller_0_s1_read                                         : out std_logic;                                        -- read
			new_sdram_controller_0_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			new_sdram_controller_0_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			new_sdram_controller_0_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			new_sdram_controller_0_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			new_sdram_controller_0_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			new_sdram_controller_0_s1_chipselect                                   : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                                   : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                                     : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                                      : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable                                : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                               : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                                            : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory2_0_s1_write                                              : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                                         : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                                         : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                                              : out std_logic;                                        -- clken
			pio_input_key_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			pio_input_key_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_input_level_s1_address                                             : out std_logic_vector(1 downto 0);                     -- address
			pio_input_level_s1_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_output_answer_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			pio_output_answer_s1_write                                             : out std_logic;                                        -- write
			pio_output_answer_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_output_answer_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			pio_output_answer_s1_chipselect                                        : out std_logic;                                        -- chipselect
			pio_sseg_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			pio_sseg_s1_write                                                      : out std_logic;                                        -- write
			pio_sseg_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_sseg_s1_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			pio_sseg_s1_chipselect                                                 : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                                     : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                                     : out std_logic_vector(2 downto 0);                     -- address
			timer_0_s1_write                                                       : out std_logic;                                        -- write
			timer_0_s1_readdata                                                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                                   : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                                  : out std_logic;                                        -- chipselect
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     : out std_logic_vector(12 downto 0);                    -- address
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       : out std_logic;                                        -- write
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        : out std_logic;                                        -- read
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  : out std_logic_vector(0 downto 0);                     -- byteenable
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  : out std_logic;                                        -- chipselect
			video_character_buffer_with_dma_0_avalon_char_control_slave_address    : out std_logic_vector(0 downto 0);                     -- address
			video_character_buffer_with_dma_0_avalon_char_control_slave_write      : out std_logic;                                        -- write
			video_character_buffer_with_dma_0_avalon_char_control_slave_read       : out std_logic;                                        -- read
			video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable : out std_logic_vector(3 downto 0);                     -- byteenable
			video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect : out std_logic                                         -- chipselect
		);
	end component finalproject_trivia_mm_interconnect_0;

	component finalproject_trivia_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component finalproject_trivia_irq_mapper;

	component finalproject_trivia_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component finalproject_trivia_rst_controller;

	component finalproject_trivia_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component finalproject_trivia_rst_controller_001;

	signal video_character_buffer_with_dma_0_avalon_char_source_valid                               : std_logic;                     -- video_character_buffer_with_dma_0:stream_valid -> video_dual_clock_buffer_0:stream_in_valid
	signal video_character_buffer_with_dma_0_avalon_char_source_data                                : std_logic_vector(29 downto 0); -- video_character_buffer_with_dma_0:stream_data -> video_dual_clock_buffer_0:stream_in_data
	signal video_character_buffer_with_dma_0_avalon_char_source_ready                               : std_logic;                     -- video_dual_clock_buffer_0:stream_in_ready -> video_character_buffer_with_dma_0:stream_ready
	signal video_character_buffer_with_dma_0_avalon_char_source_startofpacket                       : std_logic;                     -- video_character_buffer_with_dma_0:stream_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	signal video_character_buffer_with_dma_0_avalon_char_source_endofpacket                         : std_logic;                     -- video_character_buffer_with_dma_0:stream_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_valid                                  : std_logic;                     -- video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_data                                   : std_logic_vector(29 downto 0); -- video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_ready                                  : std_logic;                     -- video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket                          : std_logic;                     -- video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	signal video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket                            : std_logic;                     -- video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	signal altpll_0_c0_clk                                                                          : std_logic;                     -- altpll_0:c0 -> [irq_mapper:clk, jtag_uart_0:clk, mm_interconnect_0:altpll_0_c0_clk, new_sdram_controller_0:clk, nios2_gen2_0:clk, onchip_memory2_0:clk, rst_controller_001:clk, sysid_qsys_0:clock, timer_0:clk, video_character_buffer_with_dma_0:clk, video_dual_clock_buffer_0:clk_stream_in]
	signal altpll_0_c2_clk                                                                          : std_logic;                     -- altpll_0:c2 -> [rst_controller_002:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	signal nios2_gen2_0_data_master_readdata                                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                                     : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                                         : std_logic_vector(26 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                                      : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                                            : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                                           : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                                       : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                                              : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                                  : std_logic_vector(26 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                                     : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect -> video_character_buffer_with_dma_0:buf_chipselect
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    : std_logic_vector(7 downto 0);  -- video_character_buffer_with_dma_0:buf_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest : std_logic;                     -- video_character_buffer_with_dma_0:buf_waitrequest -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     : std_logic_vector(12 downto 0); -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_address -> video_character_buffer_with_dma_0:buf_address
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_read -> video_character_buffer_with_dma_0:buf_read
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable -> video_character_buffer_with_dma_0:buf_byteenable
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_write -> video_character_buffer_with_dma_0:buf_write
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   : std_logic_vector(7 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata -> video_character_buffer_with_dma_0:buf_writedata
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect -> video_character_buffer_with_dma_0:ctrl_chipselect
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   : std_logic_vector(31 downto 0); -- video_character_buffer_with_dma_0:ctrl_readdata -> mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_readdata
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_address -> video_character_buffer_with_dma_0:ctrl_address
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read       : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_read -> video_character_buffer_with_dma_0:ctrl_read
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable -> video_character_buffer_with_dma_0:ctrl_byteenable
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write      : std_logic;                     -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_write -> video_character_buffer_with_dma_0:ctrl_write
	signal mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_character_buffer_with_dma_0_avalon_char_control_slave_writedata -> video_character_buffer_with_dma_0:ctrl_writedata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect                               : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                                 : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest                              : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                                     : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                                    : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                                    : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                                  : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest                               : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess                               : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                                      : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable                                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                                            : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                                                : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                                               : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                                         : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                                           : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                                            : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                                         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                                              : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                                          : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                                              : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal mm_interconnect_0_timer_0_s1_chipselect                                                  : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                                                    : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                                     : std_logic_vector(2 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                                       : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                                                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_new_sdram_controller_0_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdata                                     : std_logic_vector(15 downto 0); -- new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	signal mm_interconnect_0_new_sdram_controller_0_s1_waitrequest                                  : std_logic;                     -- new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	signal mm_interconnect_0_new_sdram_controller_0_s1_address                                      : std_logic_vector(24 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	signal mm_interconnect_0_new_sdram_controller_0_s1_read                                         : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_read -> mm_interconnect_0_new_sdram_controller_0_s1_read:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> mm_interconnect_0_new_sdram_controller_0_s1_byteenable:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid                                : std_logic;                     -- new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	signal mm_interconnect_0_new_sdram_controller_0_s1_write                                        : std_logic;                     -- mm_interconnect_0:new_sdram_controller_0_s1_write -> mm_interconnect_0_new_sdram_controller_0_s1_write:in
	signal mm_interconnect_0_new_sdram_controller_0_s1_writedata                                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	signal mm_interconnect_0_pio_input_level_s1_readdata                                            : std_logic_vector(31 downto 0); -- pio_input_level:readdata -> mm_interconnect_0:pio_input_level_s1_readdata
	signal mm_interconnect_0_pio_input_level_s1_address                                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_input_level_s1_address -> pio_input_level:address
	signal mm_interconnect_0_pio_output_answer_s1_chipselect                                        : std_logic;                     -- mm_interconnect_0:pio_output_answer_s1_chipselect -> pio_output_answer:chipselect
	signal mm_interconnect_0_pio_output_answer_s1_readdata                                          : std_logic_vector(31 downto 0); -- pio_output_answer:readdata -> mm_interconnect_0:pio_output_answer_s1_readdata
	signal mm_interconnect_0_pio_output_answer_s1_address                                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_output_answer_s1_address -> pio_output_answer:address
	signal mm_interconnect_0_pio_output_answer_s1_write                                             : std_logic;                     -- mm_interconnect_0:pio_output_answer_s1_write -> mm_interconnect_0_pio_output_answer_s1_write:in
	signal mm_interconnect_0_pio_output_answer_s1_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_output_answer_s1_writedata -> pio_output_answer:writedata
	signal mm_interconnect_0_pio_input_key_s1_readdata                                              : std_logic_vector(31 downto 0); -- pio_input_key:readdata -> mm_interconnect_0:pio_input_key_s1_readdata
	signal mm_interconnect_0_pio_input_key_s1_address                                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_input_key_s1_address -> pio_input_key:address
	signal mm_interconnect_0_pio_sseg_s1_chipselect                                                 : std_logic;                     -- mm_interconnect_0:pio_sseg_s1_chipselect -> pio_sseg:chipselect
	signal mm_interconnect_0_pio_sseg_s1_readdata                                                   : std_logic_vector(31 downto 0); -- pio_sseg:readdata -> mm_interconnect_0:pio_sseg_s1_readdata
	signal mm_interconnect_0_pio_sseg_s1_address                                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_sseg_s1_address -> pio_sseg:address
	signal mm_interconnect_0_pio_sseg_s1_write                                                      : std_logic;                     -- mm_interconnect_0:pio_sseg_s1_write -> mm_interconnect_0_pio_sseg_s1_write:in
	signal mm_interconnect_0_pio_sseg_s1_writedata                                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_sseg_s1_writedata -> pio_sseg:writedata
	signal irq_mapper_receiver0_irq                                                                 : std_logic;                     -- timer_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                 : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal nios2_gen2_0_irq_irq                                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                                           : std_logic;                     -- rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset                                                       : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset, video_character_buffer_with_dma_0:reset, video_dual_clock_buffer_0:reset_stream_in]
	signal rst_controller_001_reset_out_reset_req                                                   : std_logic;                     -- rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                                                       : std_logic;                     -- rst_controller_002:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]
	signal reset_reset_n_ports_inv                                                                  : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv                           : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                                             : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv                               : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_read:inv -> new_sdram_controller_0:az_rd_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0_new_sdram_controller_0_s1_byteenable:inv -> new_sdram_controller_0:az_be_n
	signal mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_new_sdram_controller_0_s1_write:inv -> new_sdram_controller_0:az_wr_n
	signal mm_interconnect_0_pio_output_answer_s1_write_ports_inv                                   : std_logic;                     -- mm_interconnect_0_pio_output_answer_s1_write:inv -> pio_output_answer:write_n
	signal mm_interconnect_0_pio_sseg_s1_write_ports_inv                                            : std_logic;                     -- mm_interconnect_0_pio_sseg_s1_write:inv -> pio_sseg:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                 : std_logic;                     -- rst_controller_reset_out_reset:inv -> [pio_input_key:reset_n, pio_input_level:reset_n, pio_output_answer:reset_n, pio_sseg:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                             : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [jtag_uart_0:rst_n, new_sdram_controller_0:reset_n, nios2_gen2_0:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n]

begin

	altpll_0 : component finalproject_trivia_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                 -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c1                 => clk_sdram_clk,                                  --                    c1.clk
			c2                 => altpll_0_c2_clk,                                --                    c2.clk
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			c3                 => open,                                           --           (terminated)
			c4                 => open,                                           --           (terminated)
			areset             => '0',                                            --           (terminated)
			locked             => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "000",                                          --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	jtag_uart_0 : component finalproject_trivia_jtag_uart_0
		port map (
			clk            => altpll_0_c0_clk,                                                 --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                         --               irq.irq
		);

	new_sdram_controller_0 : component finalproject_trivia_new_sdram_controller_0
		port map (
			clk            => altpll_0_c0_clk,                                                  --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,                     -- reset.reset_n
			az_addr        => mm_interconnect_0_new_sdram_controller_0_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_new_sdram_controller_0_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_new_sdram_controller_0_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                                  --  wire.export
			zs_ba          => sdram_wire_ba,                                                    --      .export
			zs_cas_n       => sdram_wire_cas_n,                                                 --      .export
			zs_cke         => sdram_wire_cke,                                                   --      .export
			zs_cs_n        => sdram_wire_cs_n,                                                  --      .export
			zs_dq          => sdram_wire_dq,                                                    --      .export
			zs_dqm         => sdram_wire_dqm,                                                   --      .export
			zs_ras_n       => sdram_wire_ras_n,                                                 --      .export
			zs_we_n        => sdram_wire_we_n                                                   --      .export
		);

	nios2_gen2_0 : component finalproject_trivia_nios2_gen2_0
		port map (
			clk                                 => altpll_0_c0_clk,                                            --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,               --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,                     --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                       --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component finalproject_trivia_onchip_memory2_0
		port map (
			clk        => altpll_0_c0_clk,                                  --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,               -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,           --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	pio_input_key : component finalproject_trivia_pio_input_key
		port map (
			clk      => clk_clk,                                     --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address  => mm_interconnect_0_pio_input_key_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_input_key_s1_readdata, --                    .readdata
			in_port  => pio_input_key_external_connection_export     -- external_connection.export
		);

	pio_input_level : component finalproject_trivia_pio_input_key
		port map (
			clk      => clk_clk,                                       --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address  => mm_interconnect_0_pio_input_level_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_pio_input_level_s1_readdata, --                    .readdata
			in_port  => pio_input_level_external_connection_export     -- external_connection.export
		);

	pio_output_answer : component finalproject_trivia_pio_output_answer
		port map (
			clk        => clk_clk,                                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,               --               reset.reset_n
			address    => mm_interconnect_0_pio_output_answer_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_output_answer_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_output_answer_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_output_answer_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_output_answer_s1_readdata,        --                    .readdata
			out_port   => pio_output_answer_external_connection_export            -- external_connection.export
		);

	pio_sseg : component finalproject_trivia_pio_sseg
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_sseg_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_sseg_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_sseg_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_sseg_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_sseg_s1_readdata,        --                    .readdata
			out_port   => pio_sseg_external_connection_export            -- external_connection.export
		);

	sysid_qsys_0 : component finalproject_trivia_sysid_qsys_0
		port map (
			clock    => altpll_0_c0_clk,                                         --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,            --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component finalproject_trivia_timer_0
		port map (
			clk        => altpll_0_c0_clk,                              --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv, -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                      --   irq.irq
		);

	video_character_buffer_with_dma_0 : component finalproject_trivia_video_character_buffer_with_dma_0
		port map (
			clk                  => altpll_0_c0_clk,                                                                            --                       clk.clk
			reset                => rst_controller_001_reset_out_reset,                                                         --                     reset.reset
			ctrl_address         => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address(0),   -- avalon_char_control_slave.address
			ctrl_byteenable      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable,   --                          .byteenable
			ctrl_chipselect      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect,   --                          .chipselect
			ctrl_read            => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read,         --                          .read
			ctrl_write           => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write,        --                          .write
			ctrl_writedata       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata,    --                          .writedata
			ctrl_readdata        => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata,     --                          .readdata
			buf_byteenable       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable(0), --  avalon_char_buffer_slave.byteenable
			buf_chipselect       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect,    --                          .chipselect
			buf_read             => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read,          --                          .read
			buf_write            => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write,         --                          .write
			buf_writedata        => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata,     --                          .writedata
			buf_readdata         => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata,      --                          .readdata
			buf_waitrequest      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest,   --                          .waitrequest
			buf_address          => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address,       --                          .address
			stream_ready         => video_character_buffer_with_dma_0_avalon_char_source_ready,                                 --        avalon_char_source.ready
			stream_startofpacket => video_character_buffer_with_dma_0_avalon_char_source_startofpacket,                         --                          .startofpacket
			stream_endofpacket   => video_character_buffer_with_dma_0_avalon_char_source_endofpacket,                           --                          .endofpacket
			stream_valid         => video_character_buffer_with_dma_0_avalon_char_source_valid,                                 --                          .valid
			stream_data          => video_character_buffer_with_dma_0_avalon_char_source_data                                   --                          .data
		);

	video_dual_clock_buffer_0 : component finalproject_trivia_video_dual_clock_buffer_0
		port map (
			clk_stream_in            => altpll_0_c0_clk,                                                    --         clock_stream_in.clk
			reset_stream_in          => rst_controller_001_reset_out_reset,                                 --         reset_stream_in.reset
			clk_stream_out           => altpll_0_c2_clk,                                                    --        clock_stream_out.clk
			reset_stream_out         => rst_controller_002_reset_out_reset,                                 --        reset_stream_out.reset
			stream_in_ready          => video_character_buffer_with_dma_0_avalon_char_source_ready,         --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => video_character_buffer_with_dma_0_avalon_char_source_startofpacket, --                        .startofpacket
			stream_in_endofpacket    => video_character_buffer_with_dma_0_avalon_char_source_endofpacket,   --                        .endofpacket
			stream_in_valid          => video_character_buffer_with_dma_0_avalon_char_source_valid,         --                        .valid
			stream_in_data           => video_character_buffer_with_dma_0_avalon_char_source_data,          --                        .data
			stream_out_ready         => video_dual_clock_buffer_0_avalon_dc_buffer_source_ready,            -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket,    --                        .startofpacket
			stream_out_endofpacket   => video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,      --                        .endofpacket
			stream_out_valid         => video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,            --                        .valid
			stream_out_data          => video_dual_clock_buffer_0_avalon_dc_buffer_source_data              --                        .data
		);

	video_vga_controller_0 : component finalproject_trivia_video_vga_controller_0
		port map (
			clk           => altpll_0_c2_clk,                                                 --                clk.clk
			reset         => rst_controller_002_reset_out_reset,                              --              reset.reset
			data          => video_dual_clock_buffer_0_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => video_dual_clock_buffer_0_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => video_dual_clock_buffer_0_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_out_CLK,                                                     -- external_interface.export
			VGA_HS        => vga_out_HS,                                                      --                   .export
			VGA_VS        => vga_out_VS,                                                      --                   .export
			VGA_BLANK     => vga_out_BLANK,                                                   --                   .export
			VGA_SYNC      => vga_out_SYNC,                                                    --                   .export
			VGA_R         => vga_out_R,                                                       --                   .export
			VGA_G         => vga_out_G,                                                       --                   .export
			VGA_B         => vga_out_B                                                        --                   .export
		);

	mm_interconnect_0 : component finalproject_trivia_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                                        => altpll_0_c0_clk,                                                                          --                                                 altpll_0_c0.clk
			clk_0_clk_clk                                                          => clk_clk,                                                                                  --                                                   clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset             => rst_controller_reset_out_reset,                                                           --        altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_reset_reset_bridge_in_reset_reset                         => rst_controller_001_reset_out_reset,                                                       --                    nios2_gen2_0_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                                       => nios2_gen2_0_data_master_address,                                                         --                                    nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                                   => nios2_gen2_0_data_master_waitrequest,                                                     --                                                            .waitrequest
			nios2_gen2_0_data_master_byteenable                                    => nios2_gen2_0_data_master_byteenable,                                                      --                                                            .byteenable
			nios2_gen2_0_data_master_read                                          => nios2_gen2_0_data_master_read,                                                            --                                                            .read
			nios2_gen2_0_data_master_readdata                                      => nios2_gen2_0_data_master_readdata,                                                        --                                                            .readdata
			nios2_gen2_0_data_master_write                                         => nios2_gen2_0_data_master_write,                                                           --                                                            .write
			nios2_gen2_0_data_master_writedata                                     => nios2_gen2_0_data_master_writedata,                                                       --                                                            .writedata
			nios2_gen2_0_data_master_debugaccess                                   => nios2_gen2_0_data_master_debugaccess,                                                     --                                                            .debugaccess
			nios2_gen2_0_instruction_master_address                                => nios2_gen2_0_instruction_master_address,                                                  --                             nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest                            => nios2_gen2_0_instruction_master_waitrequest,                                              --                                                            .waitrequest
			nios2_gen2_0_instruction_master_read                                   => nios2_gen2_0_instruction_master_read,                                                     --                                                            .read
			nios2_gen2_0_instruction_master_readdata                               => nios2_gen2_0_instruction_master_readdata,                                                 --                                                            .readdata
			altpll_0_pll_slave_address                                             => mm_interconnect_0_altpll_0_pll_slave_address,                                             --                                          altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                               => mm_interconnect_0_altpll_0_pll_slave_write,                                               --                                                            .write
			altpll_0_pll_slave_read                                                => mm_interconnect_0_altpll_0_pll_slave_read,                                                --                                                            .read
			altpll_0_pll_slave_readdata                                            => mm_interconnect_0_altpll_0_pll_slave_readdata,                                            --                                                            .readdata
			altpll_0_pll_slave_writedata                                           => mm_interconnect_0_altpll_0_pll_slave_writedata,                                           --                                                            .writedata
			jtag_uart_0_avalon_jtag_slave_address                                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                                  --                               jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                                    --                                                            .write
			jtag_uart_0_avalon_jtag_slave_read                                     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                                     --                                                            .read
			jtag_uart_0_avalon_jtag_slave_readdata                                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,                                 --                                                            .readdata
			jtag_uart_0_avalon_jtag_slave_writedata                                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,                                --                                                            .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest                              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,                              --                                                            .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect                               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,                               --                                                            .chipselect
			new_sdram_controller_0_s1_address                                      => mm_interconnect_0_new_sdram_controller_0_s1_address,                                      --                                   new_sdram_controller_0_s1.address
			new_sdram_controller_0_s1_write                                        => mm_interconnect_0_new_sdram_controller_0_s1_write,                                        --                                                            .write
			new_sdram_controller_0_s1_read                                         => mm_interconnect_0_new_sdram_controller_0_s1_read,                                         --                                                            .read
			new_sdram_controller_0_s1_readdata                                     => mm_interconnect_0_new_sdram_controller_0_s1_readdata,                                     --                                                            .readdata
			new_sdram_controller_0_s1_writedata                                    => mm_interconnect_0_new_sdram_controller_0_s1_writedata,                                    --                                                            .writedata
			new_sdram_controller_0_s1_byteenable                                   => mm_interconnect_0_new_sdram_controller_0_s1_byteenable,                                   --                                                            .byteenable
			new_sdram_controller_0_s1_readdatavalid                                => mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid,                                --                                                            .readdatavalid
			new_sdram_controller_0_s1_waitrequest                                  => mm_interconnect_0_new_sdram_controller_0_s1_waitrequest,                                  --                                                            .waitrequest
			new_sdram_controller_0_s1_chipselect                                   => mm_interconnect_0_new_sdram_controller_0_s1_chipselect,                                   --                                                            .chipselect
			nios2_gen2_0_debug_mem_slave_address                                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                                   --                                nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                                     --                                                            .write
			nios2_gen2_0_debug_mem_slave_read                                      => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                                      --                                                            .read
			nios2_gen2_0_debug_mem_slave_readdata                                  => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                                  --                                                            .readdata
			nios2_gen2_0_debug_mem_slave_writedata                                 => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,                                 --                                                            .writedata
			nios2_gen2_0_debug_mem_slave_byteenable                                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,                                --                                                            .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest                               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,                               --                                                            .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess                               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,                               --                                                            .debugaccess
			onchip_memory2_0_s1_address                                            => mm_interconnect_0_onchip_memory2_0_s1_address,                                            --                                         onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                                              => mm_interconnect_0_onchip_memory2_0_s1_write,                                              --                                                            .write
			onchip_memory2_0_s1_readdata                                           => mm_interconnect_0_onchip_memory2_0_s1_readdata,                                           --                                                            .readdata
			onchip_memory2_0_s1_writedata                                          => mm_interconnect_0_onchip_memory2_0_s1_writedata,                                          --                                                            .writedata
			onchip_memory2_0_s1_byteenable                                         => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                                         --                                                            .byteenable
			onchip_memory2_0_s1_chipselect                                         => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                                         --                                                            .chipselect
			onchip_memory2_0_s1_clken                                              => mm_interconnect_0_onchip_memory2_0_s1_clken,                                              --                                                            .clken
			pio_input_key_s1_address                                               => mm_interconnect_0_pio_input_key_s1_address,                                               --                                            pio_input_key_s1.address
			pio_input_key_s1_readdata                                              => mm_interconnect_0_pio_input_key_s1_readdata,                                              --                                                            .readdata
			pio_input_level_s1_address                                             => mm_interconnect_0_pio_input_level_s1_address,                                             --                                          pio_input_level_s1.address
			pio_input_level_s1_readdata                                            => mm_interconnect_0_pio_input_level_s1_readdata,                                            --                                                            .readdata
			pio_output_answer_s1_address                                           => mm_interconnect_0_pio_output_answer_s1_address,                                           --                                        pio_output_answer_s1.address
			pio_output_answer_s1_write                                             => mm_interconnect_0_pio_output_answer_s1_write,                                             --                                                            .write
			pio_output_answer_s1_readdata                                          => mm_interconnect_0_pio_output_answer_s1_readdata,                                          --                                                            .readdata
			pio_output_answer_s1_writedata                                         => mm_interconnect_0_pio_output_answer_s1_writedata,                                         --                                                            .writedata
			pio_output_answer_s1_chipselect                                        => mm_interconnect_0_pio_output_answer_s1_chipselect,                                        --                                                            .chipselect
			pio_sseg_s1_address                                                    => mm_interconnect_0_pio_sseg_s1_address,                                                    --                                                 pio_sseg_s1.address
			pio_sseg_s1_write                                                      => mm_interconnect_0_pio_sseg_s1_write,                                                      --                                                            .write
			pio_sseg_s1_readdata                                                   => mm_interconnect_0_pio_sseg_s1_readdata,                                                   --                                                            .readdata
			pio_sseg_s1_writedata                                                  => mm_interconnect_0_pio_sseg_s1_writedata,                                                  --                                                            .writedata
			pio_sseg_s1_chipselect                                                 => mm_interconnect_0_pio_sseg_s1_chipselect,                                                 --                                                            .chipselect
			sysid_qsys_0_control_slave_address                                     => mm_interconnect_0_sysid_qsys_0_control_slave_address,                                     --                                  sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                                    => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,                                    --                                                            .readdata
			timer_0_s1_address                                                     => mm_interconnect_0_timer_0_s1_address,                                                     --                                                  timer_0_s1.address
			timer_0_s1_write                                                       => mm_interconnect_0_timer_0_s1_write,                                                       --                                                            .write
			timer_0_s1_readdata                                                    => mm_interconnect_0_timer_0_s1_readdata,                                                    --                                                            .readdata
			timer_0_s1_writedata                                                   => mm_interconnect_0_timer_0_s1_writedata,                                                   --                                                            .writedata
			timer_0_s1_chipselect                                                  => mm_interconnect_0_timer_0_s1_chipselect,                                                  --                                                            .chipselect
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_address     => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_address,     --  video_character_buffer_with_dma_0_avalon_char_buffer_slave.address
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_write       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_write,       --                                                            .write
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_read        => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_read,        --                                                            .read
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata    => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_readdata,    --                                                            .readdata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata   => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_writedata,   --                                                            .writedata
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable  => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_byteenable,  --                                                            .byteenable
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_waitrequest, --                                                            .waitrequest
			video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect  => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_buffer_slave_chipselect,  --                                                            .chipselect
			video_character_buffer_with_dma_0_avalon_char_control_slave_address    => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_address,    -- video_character_buffer_with_dma_0_avalon_char_control_slave.address
			video_character_buffer_with_dma_0_avalon_char_control_slave_write      => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_write,      --                                                            .write
			video_character_buffer_with_dma_0_avalon_char_control_slave_read       => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_read,       --                                                            .read
			video_character_buffer_with_dma_0_avalon_char_control_slave_readdata   => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_readdata,   --                                                            .readdata
			video_character_buffer_with_dma_0_avalon_char_control_slave_writedata  => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_writedata,  --                                                            .writedata
			video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_byteenable, --                                                            .byteenable
			video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect => mm_interconnect_0_video_character_buffer_with_dma_0_avalon_char_control_slave_chipselect  --                                                            .chipselect
		);

	irq_mapper : component finalproject_trivia_irq_mapper
		port map (
			clk           => altpll_0_c0_clk,                    --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq                --    sender.irq
		);

	rst_controller : component finalproject_trivia_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component finalproject_trivia_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => altpll_0_c0_clk,                        --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component finalproject_trivia_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => altpll_0_c2_clk,                    --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_new_sdram_controller_0_s1_read_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_read;

	mm_interconnect_0_new_sdram_controller_0_s1_byteenable_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_byteenable;

	mm_interconnect_0_new_sdram_controller_0_s1_write_ports_inv <= not mm_interconnect_0_new_sdram_controller_0_s1_write;

	mm_interconnect_0_pio_output_answer_s1_write_ports_inv <= not mm_interconnect_0_pio_output_answer_s1_write;

	mm_interconnect_0_pio_sseg_s1_write_ports_inv <= not mm_interconnect_0_pio_sseg_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of finalproject_trivia
